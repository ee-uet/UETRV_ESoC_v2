module user_project_wrapper (user_clock2,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    vssa2,
    vdda2,
    vssa1,
    vdda1,
    vssd2,
    vccd2,
    vssd1,
    vccd1,
    analog_io,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    user_irq,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input vssa2;
 input vdda2;
 input vssa1;
 input vdda1;
 input vssd2;
 input vccd2;
 input vssd1;
 input vccd1;
 inout [28:0] analog_io;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [127:0] la_data_in;
 output [127:0] la_data_out;
 input [127:0] la_oenb;
 output [2:0] user_irq;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;


 SoC_Tile mprj (.user_clock(user_clock2),
    .wb_clock(wb_clk_i),
    .clock_sel(io_in[5]),
    .clk_muxed(io_out[6]),
    .reset(io_in[15]),
    .io_uart_tx(io_out[29]),
    .io_uart_rx(io_in[28]),
    .io_spi_cs(io_out[26]),
    .io_spi_clk(io_out[25]),
    .io_spi_mosi(io_out[24]),
    .io_spi_miso(io_in[27]),
    .io_m1_io_qei_ch_a(io_in[7]),
    .io_m1_io_qei_ch_b(io_in[8]),
    .io_m1_io_pwm_high(io_out[9]),
    .io_m1_io_pwm_low(io_out[10]),
    .io_m1_io_x_homed(io_in[11]),
    .io_m1_io_y_homed(io_in[12]),
    .io_m1_io_step1dir(io_out[13]),
    .io_m1_io_step2dir(io_out[14]),
    .io_m2_io_qei_ch_a(io_in[16]),
    .io_m2_io_qei_ch_b(io_in[17]),
    .io_m2_io_pwm_high(io_out[18]),
    .io_m2_io_pwm_low(io_out[19]),
    .io_m2_io_x_homed(io_in[20]),
    .io_m2_io_y_homed(io_in[21]),
    .io_m2_io_step1dir(io_out[22]),
    .io_m2_io_step2dir(io_out[23]),
    .io_m3_io_qei_ch_a(io_in[30]),
    .io_m3_io_qei_ch_b(io_in[31]),
    .io_m3_io_pwm_high(io_out[32]),
    .io_m3_io_pwm_low(io_out[33]),
    .io_m3_io_x_homed(io_in[34]),
    .io_m3_io_y_homed(io_in[35]),
    .io_m3_io_step1dir(io_out[36]),
    .io_m3_io_step2dir(io_out[37]),
    .vssd1(vssd1),
    .vccd1(vccd1),
    .io_oeb({io_oeb[37],
    io_oeb[36],
    io_oeb[35],
    io_oeb[34],
    io_oeb[33],
    io_oeb[32],
    io_oeb[31],
    io_oeb[30],
    io_oeb[29],
    io_oeb[28],
    io_oeb[27],
    io_oeb[26],
    io_oeb[25],
    io_oeb[24],
    io_oeb[23],
    io_oeb[22],
    io_oeb[21],
    io_oeb[20],
    io_oeb[19],
    io_oeb[18],
    io_oeb[17],
    io_oeb[16],
    io_oeb[15],
    io_oeb[14],
    io_oeb[13],
    io_oeb[12],
    io_oeb[11],
    io_oeb[10],
    io_oeb[9],
    io_oeb[8],
    io_oeb[7],
    io_oeb[6],
    io_oeb[5],
    io_oeb[4],
    io_oeb[3],
    io_oeb[2],
    io_oeb[1],
    io_oeb[0]}));
endmodule
